class mem_mon;
	mem_tx tx;

	task run();
		$display(" #### running  run task :: MEM_MON");
		//  collect data from  interfce
		// send data to  coverage and  sbd
	endtask
endclass

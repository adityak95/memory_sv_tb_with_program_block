program mem_prgm();
mem_env env;
initial begin
	env=new();
	env.run();
end

endprogram

`define  WIDTH 8
`define  DEPTH 8
`define  ADDR_WIDTH 3
 class mem_common;
		static mailbox gen2bfm=new();
		static string  testcase="5_WRITES_5_READS";
 endclass

class mem_sbd;
	mem_tx tx;

	task run();
		$display(" #### running  run task :: MEM_SBD");
		//  collect data fro mailbox
		// compare the  tb and dut data  
	endtask
endclass

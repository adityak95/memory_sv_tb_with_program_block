class mem_cov;
	mem_tx tx;

	task run();
		$display(" #### running  run task :: MEM_COV");
		//  collect tghe dat from  mailbox
		// sample the  covergroup
	endtask
endclass
